VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ravenna
  CLASS BLOCK ;
  FOREIGN ravenna ;
  ORIGIN 0.000 0.000 ;
  SIZE 2573.000 BY 2068.000 ;
  PIN VDD3V3
    PORT
      LAYER MET1 ;
        RECT 2146.480 1962.800 2199.120 2028.880 ;
    END
  END VDD3V3
  PIN VDD1V8
    PORT
      LAYER MET1 ;
        RECT 1436.400 39.200 1489.500 104.720 ;
    END
  END VDD1V8
  PIN VSS
    PORT
      LAYER MET1 ;
        RECT 2467.880 1755.500 2533.880 1808.500 ;
    END
  END VSS
  PIN XI
    PORT
      LAYER METTPL ;
        RECT 63.840 520.800 81.200 535.920 ;
    END
  END XI
  PIN XO
    PORT
      LAYER METTPL ;
        RECT 61.600 326.480 82.320 342.720 ;
    END
  END XO
  PIN XCLK
    PORT
      LAYER MET1 ;
        RECT 2344.500 39.120 2397.500 105.120 ;
    END
  END XCLK
  PIN SDI
    PORT
      LAYER MET1 ;
        RECT 269.500 39.120 322.500 105.120 ;
    END
  END SDI
  PIN SDO
    PORT
      LAYER MET1 ;
        RECT 185.500 39.120 238.500 105.120 ;
    END
  END SDO
  PIN CSB
    PORT
      LAYER MET1 ;
        RECT 353.500 39.120 406.500 105.120 ;
    END
  END CSB
  PIN SCK
    PORT
      LAYER MET1 ;
        RECT 437.500 39.120 490.500 105.120 ;
    END
  END SCK
  PIN ser_tx
    PORT
      LAYER MET1 ;
        RECT 2467.880 1135.500 2533.880 1188.500 ;
    END
  END ser_tx
  PIN ser_rx
    PORT
      LAYER MET1 ;
        RECT 2467.880 1219.500 2533.880 1272.500 ;
    END
  END ser_rx
  PIN i2c_sda
    PORT
      LAYER MET1 ;
        RECT 2467.880 599.500 2533.880 652.500 ;
    END
  END i2c_sda
  PIN i2c_scl
    PORT
      LAYER MET1 ;
        RECT 2467.880 683.500 2533.880 736.500 ;
    END
  END i2c_scl
  PIN spi_sdi
    PORT
      LAYER MET1 ;
        RECT 2467.880 1839.500 2533.880 1892.500 ;
    END
  END spi_sdi
  PIN spi_csb
    PORT
      LAYER MET1 ;
        RECT 2467.880 1671.500 2533.880 1724.500 ;
    END
  END spi_csb
  PIN spi_sck
    PORT
      LAYER MET1 ;
        RECT 2467.880 1587.500 2533.880 1640.500 ;
    END
  END spi_sck
  PIN spi_sdo
    PORT
      LAYER MET1 ;
        RECT 2467.880 1503.500 2533.880 1556.500 ;
    END
  END spi_sdo
  PIN irq
    PORT
      LAYER MET1 ;
        RECT 2467.880 231.500 2533.880 284.500 ;
    END
  END irq
  PIN gpio[15]
    PORT
      LAYER MET1 ;
        RECT 39.200 1369.200 104.720 1422.500 ;
    END
  END gpio[15]
  PIN gpio[14]
    PORT
      LAYER MET1 ;
        RECT 39.120 1453.500 105.120 1506.500 ;
    END
  END gpio[14]
  PIN gpio[13]
    PORT
      LAYER MET1 ;
        RECT 39.120 1537.500 105.120 1590.500 ;
    END
  END gpio[13]
  PIN gpio[12]
    PORT
      LAYER MET1 ;
        RECT 39.120 1621.500 105.120 1674.500 ;
    END
  END gpio[12]
  PIN gpio[11]
    PORT
      LAYER MET1 ;
        RECT 175.840 1962.800 227.920 2028.880 ;
    END
  END gpio[11]
  PIN gpio[10]
    PORT
      LAYER MET1 ;
        RECT 259.840 1962.800 311.920 2028.880 ;
    END
  END gpio[10]
  PIN gpio[9]
    PORT
      LAYER MET1 ;
        RECT 343.840 1962.800 395.920 2028.880 ;
    END
  END gpio[9]
  PIN gpio[8]
    PORT
      LAYER MET1 ;
        RECT 427.840 1962.800 479.920 2028.880 ;
    END
  END gpio[8]
  PIN gpio[7]
    PORT
      LAYER MET1 ;
        RECT 511.840 1962.800 563.920 2028.880 ;
    END
  END gpio[7]
  PIN gpio[6]
    PORT
      LAYER MET1 ;
        RECT 595.840 1962.800 647.920 2028.880 ;
    END
  END gpio[6]
  PIN gpio[5]
    PORT
      LAYER MET1 ;
        RECT 679.840 1962.800 731.920 2028.880 ;
    END
  END gpio[5]
  PIN gpio[4]
    PORT
      LAYER MET1 ;
        RECT 963.760 1962.800 1015.840 2028.880 ;
    END
  END gpio[4]
  PIN gpio[3]
    PORT
      LAYER MET1 ;
        RECT 1047.760 1962.800 1099.840 2028.880 ;
    END
  END gpio[3]
  PIN gpio[2]
    PORT
      LAYER MET1 ;
        RECT 1182.160 1962.800 1234.240 2028.880 ;
    END
  END gpio[2]
  PIN gpio[1]
    PORT
      LAYER MET1 ;
        RECT 1266.160 1962.800 1318.240 2028.880 ;
    END
  END gpio[1]
  PIN gpio[0]
    PORT
      LAYER MET1 ;
        RECT 1349.600 1962.800 1401.680 2028.880 ;
    END
  END gpio[0]
  PIN flash_csb
    PORT
      LAYER MET1 ;
        RECT 1654.500 39.120 1707.500 105.120 ;
    END
  END flash_csb
  PIN flash_clk
    PORT
      LAYER MET1 ;
        RECT 1570.500 39.120 1623.500 105.120 ;
    END
  END flash_clk
  PIN flash_io0
    PORT
      LAYER MET1 ;
        RECT 1838.480 39.200 1891.500 104.720 ;
    END
  END flash_io0
  PIN flash_io1
    PORT
      LAYER MET1 ;
        RECT 1922.480 39.200 1975.500 104.720 ;
    END
  END flash_io1
  PIN flash_io2
    PORT
      LAYER MET1 ;
        RECT 2006.480 39.200 2059.500 104.720 ;
    END
  END flash_io2
  PIN flash_io3
    PORT
      LAYER MET1 ;
        RECT 2090.480 39.200 2143.500 104.720 ;
    END
  END flash_io3
  PIN adc_high
    PORT
      LAYER MET1 ;
        RECT 39.120 971.500 105.120 1024.500 ;
    END
  END adc_high
  PIN adc_low
    PORT
      LAYER MET1 ;
        RECT 39.120 887.500 105.120 940.500 ;
    END
  END adc_low
  PIN adc0_in
    PORT
      LAYER MET1 ;
        RECT 39.120 719.500 105.120 772.500 ;
    END
  END adc0_in
  PIN adc1_in
    PORT
      LAYER MET1 ;
        RECT 39.120 803.500 105.120 856.500 ;
    END
  END adc1_in
  PIN analog_out
    PORT
      LAYER MET1 ;
        RECT 39.120 1055.500 105.120 1108.500 ;
    END
  END analog_out
  PIN comp_inp
    PORT
      LAYER MET1 ;
        RECT 39.120 1223.500 105.120 1276.500 ;
    END
  END comp_inp
  PIN comp_inn
    PORT
      LAYER MET1 ;
        RECT 39.120 1139.500 105.120 1192.500 ;
    END
  END comp_inn
  PIN nvref_ext
    PORT
      LAYER MET1 ;
        RECT 39.120 585.500 105.120 638.500 ;
    END
  END nvref_ext
  OBS
      LAYER MET1 ;
        RECT 0.000 2029.480 2573.000 2068.000 ;
        RECT 0.000 1962.200 175.240 2029.480 ;
        RECT 228.520 1962.200 259.240 2029.480 ;
        RECT 312.520 1962.200 343.240 2029.480 ;
        RECT 396.520 1962.200 427.240 2029.480 ;
        RECT 480.520 1962.200 511.240 2029.480 ;
        RECT 564.520 1962.200 595.240 2029.480 ;
        RECT 648.520 1962.200 679.240 2029.480 ;
        RECT 732.520 1962.200 963.160 2029.480 ;
        RECT 1016.440 1962.200 1047.160 2029.480 ;
        RECT 1100.440 1962.200 1181.560 2029.480 ;
        RECT 1234.840 1962.200 1265.560 2029.480 ;
        RECT 1318.840 1962.200 1349.000 2029.480 ;
        RECT 1402.280 1962.200 2145.880 2029.480 ;
        RECT 2199.720 1962.200 2573.000 2029.480 ;
        RECT 0.000 1893.100 2573.000 1962.200 ;
        RECT 0.000 1838.900 2467.280 1893.100 ;
        RECT 2534.480 1838.900 2573.000 1893.100 ;
        RECT 0.000 1809.100 2573.000 1838.900 ;
        RECT 0.000 1754.900 2467.280 1809.100 ;
        RECT 2534.480 1754.900 2573.000 1809.100 ;
        RECT 0.000 1725.100 2573.000 1754.900 ;
        RECT 0.000 1675.100 2467.280 1725.100 ;
        RECT 0.000 1620.900 38.520 1675.100 ;
        RECT 105.720 1670.900 2467.280 1675.100 ;
        RECT 2534.480 1670.900 2573.000 1725.100 ;
        RECT 105.720 1641.100 2573.000 1670.900 ;
        RECT 105.720 1620.900 2467.280 1641.100 ;
        RECT 0.000 1591.100 2467.280 1620.900 ;
        RECT 0.000 1536.900 38.520 1591.100 ;
        RECT 105.720 1586.900 2467.280 1591.100 ;
        RECT 2534.480 1586.900 2573.000 1641.100 ;
        RECT 105.720 1557.100 2573.000 1586.900 ;
        RECT 105.720 1536.900 2467.280 1557.100 ;
        RECT 0.000 1507.100 2467.280 1536.900 ;
        RECT 0.000 1452.900 38.520 1507.100 ;
        RECT 105.720 1502.900 2467.280 1507.100 ;
        RECT 2534.480 1502.900 2573.000 1557.100 ;
        RECT 105.720 1452.900 2573.000 1502.900 ;
        RECT 0.000 1423.100 2573.000 1452.900 ;
        RECT 0.000 1368.600 38.600 1423.100 ;
        RECT 105.320 1368.600 2573.000 1423.100 ;
        RECT 0.000 1277.100 2573.000 1368.600 ;
        RECT 0.000 1222.900 38.520 1277.100 ;
        RECT 105.720 1273.100 2573.000 1277.100 ;
        RECT 105.720 1222.900 2467.280 1273.100 ;
        RECT 0.000 1218.900 2467.280 1222.900 ;
        RECT 2534.480 1218.900 2573.000 1273.100 ;
        RECT 0.000 1193.100 2573.000 1218.900 ;
        RECT 0.000 1138.900 38.520 1193.100 ;
        RECT 105.720 1189.100 2573.000 1193.100 ;
        RECT 105.720 1138.900 2467.280 1189.100 ;
        RECT 0.000 1134.900 2467.280 1138.900 ;
        RECT 2534.480 1134.900 2573.000 1189.100 ;
        RECT 0.000 1109.100 2573.000 1134.900 ;
        RECT 0.000 1054.900 38.520 1109.100 ;
        RECT 105.720 1054.900 2573.000 1109.100 ;
        RECT 0.000 1025.100 2573.000 1054.900 ;
        RECT 0.000 970.900 38.520 1025.100 ;
        RECT 105.720 970.900 2573.000 1025.100 ;
        RECT 0.000 941.100 2573.000 970.900 ;
        RECT 0.000 886.900 38.520 941.100 ;
        RECT 105.720 886.900 2573.000 941.100 ;
        RECT 0.000 857.100 2573.000 886.900 ;
        RECT 0.000 802.900 38.520 857.100 ;
        RECT 105.720 802.900 2573.000 857.100 ;
        RECT 0.000 773.100 2573.000 802.900 ;
        RECT 0.000 718.900 38.520 773.100 ;
        RECT 105.720 737.100 2573.000 773.100 ;
        RECT 105.720 718.900 2467.280 737.100 ;
        RECT 0.000 682.900 2467.280 718.900 ;
        RECT 2534.480 682.900 2573.000 737.100 ;
        RECT 0.000 653.100 2573.000 682.900 ;
        RECT 0.000 639.100 2467.280 653.100 ;
        RECT 0.000 584.900 38.520 639.100 ;
        RECT 105.720 598.900 2467.280 639.100 ;
        RECT 2534.480 598.900 2573.000 653.100 ;
        RECT 105.720 584.900 2573.000 598.900 ;
        RECT 0.000 285.100 2573.000 584.900 ;
        RECT 0.000 230.900 2467.280 285.100 ;
        RECT 2534.480 230.900 2573.000 285.100 ;
        RECT 0.000 105.720 2573.000 230.900 ;
        RECT 0.000 38.520 184.900 105.720 ;
        RECT 239.100 38.520 268.900 105.720 ;
        RECT 323.100 38.520 352.900 105.720 ;
        RECT 407.100 38.520 436.900 105.720 ;
        RECT 491.100 105.320 1569.900 105.720 ;
        RECT 491.100 38.600 1435.800 105.320 ;
        RECT 1490.100 38.600 1569.900 105.320 ;
        RECT 491.100 38.520 1569.900 38.600 ;
        RECT 1624.100 38.520 1653.900 105.720 ;
        RECT 1708.100 105.320 2343.900 105.720 ;
        RECT 1708.100 38.600 1837.880 105.320 ;
        RECT 1892.100 38.600 1921.880 105.320 ;
        RECT 1976.100 38.600 2005.880 105.320 ;
        RECT 2060.100 38.600 2089.880 105.320 ;
        RECT 2144.100 38.600 2343.900 105.320 ;
        RECT 1708.100 38.520 2343.900 38.600 ;
        RECT 2398.100 38.520 2573.000 105.720 ;
        RECT 0.000 0.000 2573.000 38.520 ;
      LAYER MET2 ;
        RECT 0.000 0.000 2573.000 2068.000 ;
      LAYER MET3 ;
        RECT 0.000 0.000 2573.000 2068.000 ;
      LAYER MET4 ;
        RECT 0.000 0.000 2573.000 2068.000 ;
      LAYER METTP ;
        RECT 0.000 0.000 2573.000 2068.000 ;
      LAYER METTPL ;
        RECT 0.000 538.420 2573.000 2068.000 ;
        RECT 0.000 518.300 61.340 538.420 ;
        RECT 83.700 518.300 2573.000 538.420 ;
        RECT 0.000 345.220 2573.000 518.300 ;
        RECT 0.000 323.980 59.100 345.220 ;
        RECT 84.820 323.980 2573.000 345.220 ;
        RECT 0.000 0.000 2573.000 323.980 ;
  END
END ravenna
END LIBRARY

