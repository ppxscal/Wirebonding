VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

MACRO frequency_divid
  CLASS BLOCK ;
  FOREIGN frequency_divid ;
  ORIGIN 0.000 0.000 ;
  SIZE 664.000 BY 664.000 ;
  PIN RESET
    PORT
      LAYER met5 ;
        RECT 32.990 220.200 95.440 282.800 ;
    END
  END RESET
  PIN IN
    PORT
      LAYER met5 ;
        RECT 32.990 305.200 95.440 367.800 ;
    END
  END IN
  PIN OUT
    PORT
      LAYER met5 ;
        RECT 32.990 390.200 95.440 452.800 ;
    END
  END OUT
  PIN VDD3V3
    PORT
      LAYER met5 ;
        RECT 218.100 568.010 280.800 630.625 ;
    END
  END VDD3V3
  PIN VDD1V8
    PORT
      LAYER met5 ;
        RECT 302.100 568.010 364.800 630.625 ;
    END
  END VDD1V8
  PIN GND
    PORT
      LAYER met5 ;
        RECT 386.100 568.010 448.800 630.625 ;
    END
  END GND
  PIN N[0]
    PORT
      LAYER met5 ;
        RECT 568.560 381.200 631.010 443.800 ;
    END
  END N[0]
  PIN N[1]
    PORT
      LAYER met5 ;
        RECT 568.560 296.200 631.010 358.800 ;
    END
  END N[1]
  PIN N[2]
    PORT
      LAYER met5 ;
        RECT 568.560 211.200 631.010 273.800 ;
    END
  END N[2]
  PIN N[3]
    PORT
      LAYER met5 ;
        RECT 381.200 32.990 443.800 95.440 ;
    END
  END N[3]
  PIN N[4]
    PORT
      LAYER met5 ;
        RECT 296.200 32.990 358.800 95.440 ;
    END
  END N[4]
  PIN N[5]
    PORT
      LAYER met5 ;
        RECT 211.200 32.990 273.800 95.440 ;
    END
  END N[5]
  OBS
      LAYER li1 ;
        RECT 0.295 0.295 663.705 663.695 ;
      LAYER met1 ;
        RECT 0.000 0.000 664.000 663.725 ;
      LAYER met2 ;
        RECT 0.000 0.000 664.000 659.075 ;
      LAYER met3 ;
        RECT 0.000 0.000 664.000 664.000 ;
      LAYER met4 ;
        RECT 0.000 0.000 664.000 664.000 ;
      LAYER met5 ;
        RECT 0.000 632.225 664.000 664.000 ;
        RECT 0.000 566.410 216.500 632.225 ;
        RECT 282.400 566.410 300.500 632.225 ;
        RECT 366.400 566.410 384.500 632.225 ;
        RECT 450.400 566.410 664.000 632.225 ;
        RECT 0.000 454.400 664.000 566.410 ;
        RECT 0.000 388.600 31.390 454.400 ;
        RECT 97.040 445.400 664.000 454.400 ;
        RECT 97.040 388.600 566.960 445.400 ;
        RECT 0.000 379.600 566.960 388.600 ;
        RECT 632.610 379.600 664.000 445.400 ;
        RECT 0.000 369.400 664.000 379.600 ;
        RECT 0.000 303.600 31.390 369.400 ;
        RECT 97.040 360.400 664.000 369.400 ;
        RECT 97.040 303.600 566.960 360.400 ;
        RECT 0.000 294.600 566.960 303.600 ;
        RECT 632.610 294.600 664.000 360.400 ;
        RECT 0.000 284.400 664.000 294.600 ;
        RECT 0.000 218.600 31.390 284.400 ;
        RECT 97.040 275.400 664.000 284.400 ;
        RECT 97.040 218.600 566.960 275.400 ;
        RECT 0.000 209.600 566.960 218.600 ;
        RECT 632.610 209.600 664.000 275.400 ;
        RECT 0.000 97.040 664.000 209.600 ;
        RECT 0.000 31.390 209.600 97.040 ;
        RECT 275.400 31.390 294.600 97.040 ;
        RECT 360.400 31.390 379.600 97.040 ;
        RECT 445.400 31.390 664.000 97.040 ;
        RECT 0.000 0.000 664.000 31.390 ;
  END
END frequency_divid
