VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO raven
  CLASS BLOCK ;
  FOREIGN raven ;
  ORIGIN 608.650 97.260 ;
  SIZE 1939.000 BY 1699.000 ;
  PIN VDD3V3
    PORT
      LAYER MET1 ;
        RECT 1225.230 652.240 1291.230 705.240 ;
    END
  END VDD3V3
  PIN VDD1V8
    PORT
      LAYER MET1 ;
        RECT 1225.230 736.240 1291.230 789.240 ;
    END
  END VDD1V8
  PIN VSS
    PORT
      LAYER MET1 ;
        RECT 1225.230 568.240 1291.230 621.240 ;
    END
  END VSS
  PIN XCLK
    PORT
      LAYER MET1 ;
        RECT 768.850 -58.140 821.850 7.860 ;
    END
  END XCLK
  PIN SDI
    PORT
      LAYER MET1 ;
        RECT -220.150 -58.140 -167.150 7.860 ;
    END
  END SDI
  PIN SDO
    PORT
      LAYER MET1 ;
        RECT 51.850 -58.140 104.850 7.860 ;
    END
  END SDO
  PIN CSB
    PORT
      LAYER MET1 ;
        RECT -116.150 -58.140 -63.150 7.860 ;
    END
  END CSB
  PIN SCK
    PORT
      LAYER MET1 ;
        RECT -32.150 -58.140 20.850 7.860 ;
    END
  END SCK
  PIN ser_tx
    PORT
      LAYER MET1 ;
        RECT 1225.230 182.240 1291.230 235.240 ;
    END
  END ser_tx
  PIN ser_rx
    PORT
      LAYER MET1 ;
        RECT 1225.230 98.240 1291.230 151.240 ;
    END
  END ser_rx
  PIN irq
    PORT
      LAYER MET1 ;
        RECT 1225.230 266.240 1291.230 319.240 ;
    END
  END irq
  PIN gpio[15]
    PORT
      LAYER MET1 ;
        RECT -329.150 -58.140 -276.150 7.860 ;
    END
  END gpio[15]
  PIN gpio[14]
    PORT
      LAYER MET1 ;
        RECT -569.530 247.240 -503.530 300.240 ;
    END
  END gpio[14]
  PIN gpio[13]
    PORT
      LAYER MET1 ;
        RECT -569.530 331.240 -503.530 384.240 ;
    END
  END gpio[13]
  PIN gpio[12]
    PORT
      LAYER MET1 ;
        RECT -569.530 415.240 -503.530 468.240 ;
    END
  END gpio[12]
  PIN gpio[11]
    PORT
      LAYER MET1 ;
        RECT -569.530 499.240 -503.530 552.240 ;
    END
  END gpio[11]
  PIN gpio[10]
    PORT
      LAYER MET1 ;
        RECT -569.530 583.240 -503.530 636.240 ;
    END
  END gpio[10]
  PIN gpio[9]
    PORT
      LAYER MET1 ;
        RECT -569.530 667.240 -503.530 720.240 ;
    END
  END gpio[9]
  PIN gpio[8]
    PORT
      LAYER MET1 ;
        RECT -569.530 751.240 -503.530 804.240 ;
    END
  END gpio[8]
  PIN gpio[7]
    PORT
      LAYER MET1 ;
        RECT -569.530 835.240 -503.530 888.240 ;
    END
  END gpio[7]
  PIN gpio[6]
    PORT
      LAYER MET1 ;
        RECT -569.530 919.240 -503.530 972.240 ;
    END
  END gpio[6]
  PIN gpio[5]
    PORT
      LAYER MET1 ;
        RECT -569.530 1003.240 -503.530 1056.240 ;
    END
  END gpio[5]
  PIN gpio[4]
    PORT
      LAYER MET1 ;
        RECT -569.530 1087.240 -503.530 1140.240 ;
    END
  END gpio[4]
  PIN gpio[3]
    PORT
      LAYER MET1 ;
        RECT -569.530 1171.240 -503.530 1224.240 ;
    END
  END gpio[3]
  PIN gpio[2]
    PORT
      LAYER MET1 ;
        RECT -413.150 1496.620 -360.150 1562.620 ;
    END
  END gpio[2]
  PIN gpio[1]
    PORT
      LAYER MET1 ;
        RECT -329.150 1496.620 -276.150 1562.620 ;
    END
  END gpio[1]
  PIN gpio[0]
    PORT
      LAYER MET1 ;
        RECT -245.150 1496.620 -192.150 1562.620 ;
    END
  END gpio[0]
  PIN flash_csb
    PORT
      LAYER MET1 ;
        RECT 600.850 -58.140 653.850 7.860 ;
    END
  END flash_csb
  PIN flash_clk
    PORT
      LAYER MET1 ;
        RECT 684.850 -58.140 737.850 7.860 ;
    END
  END flash_clk
  PIN flash_io0
    PORT
      LAYER MET1 ;
        RECT 516.850 -58.140 569.850 7.860 ;
    END
  END flash_io0
  PIN flash_io1
    PORT
      LAYER MET1 ;
        RECT 432.850 -58.140 485.850 7.860 ;
    END
  END flash_io1
  PIN flash_io2
    PORT
      LAYER MET1 ;
        RECT 348.850 -58.140 401.850 7.860 ;
    END
  END flash_io2
  PIN flash_io3
    PORT
      LAYER MET1 ;
        RECT 264.850 -58.140 317.850 7.860 ;
    END
  END flash_io3
  PIN adc_high
    PORT
      LAYER MET1 ;
        RECT 997.850 1496.620 1050.850 1562.620 ;
    END
  END adc_high
  PIN adc_low
    PORT
      LAYER MET1 ;
        RECT 913.850 1496.620 966.850 1562.620 ;
    END
  END adc_low
  PIN adc0_in
    PORT
      LAYER MET1 ;
        RECT 745.850 1496.620 798.850 1562.620 ;
    END
  END adc0_in
  PIN adc1_in
    PORT
      LAYER MET1 ;
        RECT 829.850 1496.620 882.850 1562.620 ;
    END
  END adc1_in
  PIN analog_out
    PORT
      LAYER MET1 ;
        RECT 1081.850 1496.620 1134.850 1562.620 ;
    END
  END analog_out
  PIN comp_inp
    PORT
      LAYER MET1 ;
        RECT 1225.230 350.240 1291.230 403.240 ;
    END
  END comp_inp
  PIN comp_inn
    PORT
      LAYER MET1 ;
        RECT 1225.230 434.240 1291.230 487.240 ;
    END
  END comp_inn
  PIN XI
    PORT
      LAYER METTPL ;
        RECT 50.145 1521.230 64.680 1537.655 ;
    END
  END XI
  PIN XO
    PORT
      LAYER METTPL ;
        RECT -143.330 1522.330 -128.550 1538.590 ;
    END
  END XO
  OBS
      LAYER MET1 ;
        RECT -608.650 1563.220 1330.350 1601.740 ;
        RECT -608.650 1496.020 -413.750 1563.220 ;
        RECT -359.550 1496.020 -329.750 1563.220 ;
        RECT -275.550 1496.020 -245.750 1563.220 ;
        RECT -191.550 1496.020 745.250 1563.220 ;
        RECT 799.450 1496.020 829.250 1563.220 ;
        RECT 883.450 1496.020 913.250 1563.220 ;
        RECT 967.450 1496.020 997.250 1563.220 ;
        RECT 1051.450 1496.020 1081.250 1563.220 ;
        RECT 1135.450 1496.020 1330.350 1563.220 ;
        RECT -608.650 1224.840 1330.350 1496.020 ;
        RECT -608.650 1170.640 -570.130 1224.840 ;
        RECT -502.930 1170.640 1330.350 1224.840 ;
        RECT -608.650 1140.840 1330.350 1170.640 ;
        RECT -608.650 1086.640 -570.130 1140.840 ;
        RECT -502.930 1086.640 1330.350 1140.840 ;
        RECT -608.650 1056.840 1330.350 1086.640 ;
        RECT -608.650 1002.640 -570.130 1056.840 ;
        RECT -502.930 1002.640 1330.350 1056.840 ;
        RECT -608.650 972.840 1330.350 1002.640 ;
        RECT -608.650 918.640 -570.130 972.840 ;
        RECT -502.930 918.640 1330.350 972.840 ;
        RECT -608.650 888.840 1330.350 918.640 ;
        RECT -608.650 834.640 -570.130 888.840 ;
        RECT -502.930 834.640 1330.350 888.840 ;
        RECT -608.650 804.840 1330.350 834.640 ;
        RECT -608.650 750.640 -570.130 804.840 ;
        RECT -502.930 789.840 1330.350 804.840 ;
        RECT -502.930 750.640 1224.630 789.840 ;
        RECT -608.650 735.640 1224.630 750.640 ;
        RECT 1291.830 735.640 1330.350 789.840 ;
        RECT -608.650 720.840 1330.350 735.640 ;
        RECT -608.650 666.640 -570.130 720.840 ;
        RECT -502.930 705.840 1330.350 720.840 ;
        RECT -502.930 666.640 1224.630 705.840 ;
        RECT -608.650 651.640 1224.630 666.640 ;
        RECT 1291.830 651.640 1330.350 705.840 ;
        RECT -608.650 636.840 1330.350 651.640 ;
        RECT -608.650 582.640 -570.130 636.840 ;
        RECT -502.930 621.840 1330.350 636.840 ;
        RECT -502.930 582.640 1224.630 621.840 ;
        RECT -608.650 567.640 1224.630 582.640 ;
        RECT 1291.830 567.640 1330.350 621.840 ;
        RECT -608.650 552.840 1330.350 567.640 ;
        RECT -608.650 498.640 -570.130 552.840 ;
        RECT -502.930 498.640 1330.350 552.840 ;
        RECT -608.650 487.840 1330.350 498.640 ;
        RECT -608.650 468.840 1224.630 487.840 ;
        RECT -608.650 414.640 -570.130 468.840 ;
        RECT -502.930 433.640 1224.630 468.840 ;
        RECT 1291.830 433.640 1330.350 487.840 ;
        RECT -502.930 414.640 1330.350 433.640 ;
        RECT -608.650 403.840 1330.350 414.640 ;
        RECT -608.650 384.840 1224.630 403.840 ;
        RECT -608.650 330.640 -570.130 384.840 ;
        RECT -502.930 349.640 1224.630 384.840 ;
        RECT 1291.830 349.640 1330.350 403.840 ;
        RECT -502.930 330.640 1330.350 349.640 ;
        RECT -608.650 319.840 1330.350 330.640 ;
        RECT -608.650 300.840 1224.630 319.840 ;
        RECT -608.650 246.640 -570.130 300.840 ;
        RECT -502.930 265.640 1224.630 300.840 ;
        RECT 1291.830 265.640 1330.350 319.840 ;
        RECT -502.930 246.640 1330.350 265.640 ;
        RECT -608.650 235.840 1330.350 246.640 ;
        RECT -608.650 181.640 1224.630 235.840 ;
        RECT 1291.830 181.640 1330.350 235.840 ;
        RECT -608.650 151.840 1330.350 181.640 ;
        RECT -608.650 97.640 1224.630 151.840 ;
        RECT 1291.830 97.640 1330.350 151.840 ;
        RECT -608.650 8.460 1330.350 97.640 ;
        RECT -608.650 -58.740 -329.750 8.460 ;
        RECT -275.550 -58.740 -220.750 8.460 ;
        RECT -166.550 -58.740 -116.750 8.460 ;
        RECT -62.550 -58.740 -32.750 8.460 ;
        RECT 21.450 -58.740 51.250 8.460 ;
        RECT 105.450 -58.740 264.250 8.460 ;
        RECT 318.450 -58.740 348.250 8.460 ;
        RECT 402.450 -58.740 432.250 8.460 ;
        RECT 486.450 -58.740 516.250 8.460 ;
        RECT 570.450 -58.740 600.250 8.460 ;
        RECT 654.450 -58.740 684.250 8.460 ;
        RECT 738.450 -58.740 768.250 8.460 ;
        RECT 822.450 -58.740 1330.350 8.460 ;
        RECT -608.650 -97.260 1330.350 -58.740 ;
      LAYER MET2 ;
        RECT -608.650 -97.260 1330.350 1601.740 ;
      LAYER MET3 ;
        RECT -608.650 -97.260 1330.350 1601.740 ;
      LAYER MET4 ;
        RECT -608.650 -97.260 1330.350 1601.740 ;
      LAYER METTP ;
        RECT -608.650 -97.260 1330.350 1601.740 ;
      LAYER METTPL ;
        RECT -608.650 1541.090 1330.350 1601.740 ;
        RECT -608.650 1519.830 -145.830 1541.090 ;
        RECT -126.050 1540.155 1330.350 1541.090 ;
        RECT -126.050 1519.830 47.645 1540.155 ;
        RECT -608.650 1518.730 47.645 1519.830 ;
        RECT 67.180 1518.730 1330.350 1540.155 ;
        RECT -608.650 -97.260 1330.350 1518.730 ;
  END
END raven
END LIBRARY

