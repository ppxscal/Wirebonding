VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO openram_tc_1kb
  CLASS BLOCK ;
  FOREIGN openram_tc_1kb ;
  ORIGIN 0.000 0.000 ;
  SIZE 4430.000 BY 4945.000 ;
  PIN clk0
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 1240.200 3577.060 1302.800 3639.510 ;
    END
  END clk0
  PIN addr0[0]
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 1330.200 3577.060 1392.800 3639.510 ;
    END
  END addr0[0]
  PIN wmask0[3]
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 1420.200 3577.060 1482.800 3639.510 ;
    END
  END wmask0[3]
  PIN wmask0[2]
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 1511.200 3577.060 1573.800 3639.510 ;
    END
  END wmask0[2]
  PIN wmask0[1]
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 1601.200 3577.060 1663.800 3639.510 ;
    END
  END wmask0[1]
  PIN wmask0[0]
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 1691.200 3577.060 1753.800 3639.510 ;
    END
  END wmask0[0]
  PIN din0_0
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 1781.200 3577.060 1843.800 3639.510 ;
    END
  END din0_0
  PIN dout0_0
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met5 ;
        RECT 1872.200 3577.060 1934.800 3639.510 ;
    END
  END dout0_0
  PIN dout0_7
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met5 ;
        RECT 1962.200 3577.060 2024.800 3639.510 ;
    END
  END dout0_7
  PIN din0_7
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 2052.200 3577.060 2114.800 3639.510 ;
    END
  END din0_7
  PIN dout0_8
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met5 ;
        RECT 2142.200 3577.060 2204.800 3639.510 ;
    END
  END dout0_8
  PIN din0_8
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 2233.200 3577.060 2295.800 3639.510 ;
    END
  END din0_8
  PIN din0_15
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 2323.200 3577.060 2385.800 3639.510 ;
    END
  END din0_15
  PIN dout0_15
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met5 ;
        RECT 2413.200 3577.060 2475.800 3639.510 ;
    END
  END dout0_15
  PIN din0_16
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 2503.200 3577.060 2565.800 3639.510 ;
    END
  END din0_16
  PIN dout0_16
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met5 ;
        RECT 2594.200 3577.060 2656.800 3639.510 ;
    END
  END dout0_16
  PIN din0_23
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 2684.200 3577.060 2746.800 3639.510 ;
    END
  END din0_23
  PIN dout0_23
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met5 ;
        RECT 2774.200 3577.060 2836.800 3639.510 ;
    END
  END dout0_23
  PIN din0_24
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 2864.200 3577.060 2926.800 3639.510 ;
    END
  END din0_24
  PIN dout0_24
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met5 ;
        RECT 2955.200 3577.060 3017.800 3639.510 ;
    END
  END dout0_24
  PIN din0_31
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 3045.200 3577.060 3107.800 3639.510 ;
    END
  END din0_31
  PIN dout0_31
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met5 ;
        RECT 3135.200 3577.060 3197.800 3639.510 ;
    END
  END dout0_31
  PIN dout1_8
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met5 ;
        RECT 1258.200 1305.490 1320.800 1367.940 ;
    END
  END dout1_8
  PIN dout1_7
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met5 ;
        RECT 1375.200 1305.490 1437.800 1367.940 ;
    END
  END dout1_7
  PIN dout1_31
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met5 ;
        RECT 1492.200 1305.490 1554.800 1367.940 ;
    END
  END dout1_31
  PIN dout1_24
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met5 ;
        RECT 1610.200 1305.490 1672.800 1367.940 ;
    END
  END dout1_24
  PIN dout1_23
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met5 ;
        RECT 1727.200 1305.490 1789.800 1367.940 ;
    END
  END dout1_23
  PIN dout1_16
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met5 ;
        RECT 1844.200 1305.490 1906.800 1367.940 ;
    END
  END dout1_16
  PIN dout1_15
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met5 ;
        RECT 1961.200 1305.490 2023.800 1367.940 ;
    END
  END dout1_15
  PIN dout1_0
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met5 ;
        RECT 2079.200 1305.490 2141.800 1367.940 ;
    END
  END dout1_0
  PIN addr1[0]
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 2196.200 1305.490 2258.800 1367.940 ;
    END
  END addr1[0]
  PIN clk1
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 2313.200 1305.490 2375.800 1367.940 ;
    END
  END clk1
  PIN vdd
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT 2655.200 1305.875 2717.900 1368.490 ;
    END
  END vdd
  PIN vdd1v8
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT 3104.200 1305.875 3166.900 1368.490 ;
    END
  END vdd1v8
  PIN addr0[7]
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 1047.990 1547.700 1110.440 1610.300 ;
    END
  END addr0[7]
  PIN addr0[6]
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 1047.990 1687.700 1110.440 1750.300 ;
    END
  END addr0[6]
  PIN addr0[5]
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 1047.990 1827.700 1110.440 1890.300 ;
    END
  END addr0[5]
  PIN addr0[4]
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 1047.990 1967.700 1110.440 2030.300 ;
    END
  END addr0[4]
  PIN addr0[3]
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 1047.990 2107.700 1110.440 2170.300 ;
    END
  END addr0[3]
  PIN addr0[2]
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 1047.990 2247.700 1110.440 2310.300 ;
    END
  END addr0[2]
  PIN addr0[1]
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 1047.990 2387.700 1110.440 2450.300 ;
    END
  END addr0[1]
  PIN web0
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 1047.990 2527.700 1110.440 2590.300 ;
    END
  END web0
  PIN csb0
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 1047.990 2667.700 1110.440 2730.300 ;
    END
  END csb0
  PIN vss
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT 1048.375 2802.600 1110.990 2865.300 ;
    END
  END vss
  PIN csb1
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 3319.560 1529.700 3382.010 1592.300 ;
    END
  END csb1
  PIN addr1[1]
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 3319.560 1661.700 3382.010 1724.300 ;
    END
  END addr1[1]
  PIN addr1[2]
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 3319.560 1793.700 3382.010 1856.300 ;
    END
  END addr1[2]
  PIN addr1[3]
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 3319.560 1925.700 3382.010 1988.300 ;
    END
  END addr1[3]
  PIN addr1[4]
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 3319.560 2057.700 3382.010 2120.300 ;
    END
  END addr1[4]
  PIN addr1[5]
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 3319.560 2189.700 3382.010 2252.300 ;
    END
  END addr1[5]
  PIN addr1[6]
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 3319.560 2321.700 3382.010 2384.300 ;
    END
  END addr1[6]
  PIN addr1[7]
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 3319.560 2453.700 3382.010 2516.300 ;
    END
  END addr1[7]
  OBS
      LAYER li1 ;
        RECT 1.000 1.000 4429.000 4944.000 ;
      LAYER met1 ;
        RECT 1.800 1.800 4428.200 4943.200 ;
      LAYER met2 ;
        RECT 1015.000 1272.500 3415.000 3672.500 ;
      LAYER met3 ;
        RECT 1015.000 1272.500 3415.000 3672.500 ;
      LAYER met4 ;
        RECT 1015.000 1272.500 3415.000 3672.500 ;
      LAYER met5 ;
        RECT 1015.000 3641.110 3415.000 3672.500 ;
        RECT 1015.000 3575.460 1238.600 3641.110 ;
        RECT 1304.400 3575.460 1328.600 3641.110 ;
        RECT 1394.400 3575.460 1418.600 3641.110 ;
        RECT 1484.400 3575.460 1509.600 3641.110 ;
        RECT 1575.400 3575.460 1599.600 3641.110 ;
        RECT 1665.400 3575.460 1689.600 3641.110 ;
        RECT 1755.400 3575.460 1779.600 3641.110 ;
        RECT 1845.400 3575.460 1870.600 3641.110 ;
        RECT 1936.400 3575.460 1960.600 3641.110 ;
        RECT 2026.400 3575.460 2050.600 3641.110 ;
        RECT 2116.400 3575.460 2140.600 3641.110 ;
        RECT 2206.400 3575.460 2231.600 3641.110 ;
        RECT 2297.400 3575.460 2321.600 3641.110 ;
        RECT 2387.400 3575.460 2411.600 3641.110 ;
        RECT 2477.400 3575.460 2501.600 3641.110 ;
        RECT 2567.400 3575.460 2592.600 3641.110 ;
        RECT 2658.400 3575.460 2682.600 3641.110 ;
        RECT 2748.400 3575.460 2772.600 3641.110 ;
        RECT 2838.400 3575.460 2862.600 3641.110 ;
        RECT 2928.400 3575.460 2953.600 3641.110 ;
        RECT 3019.400 3575.460 3043.600 3641.110 ;
        RECT 3109.400 3575.460 3133.600 3641.110 ;
        RECT 3199.400 3575.460 3415.000 3641.110 ;
        RECT 1015.000 2866.900 3415.000 3575.460 ;
        RECT 1015.000 2801.000 1046.775 2866.900 ;
        RECT 1112.590 2801.000 3415.000 2866.900 ;
        RECT 1015.000 2731.900 3415.000 2801.000 ;
        RECT 1015.000 2666.100 1046.390 2731.900 ;
        RECT 1112.040 2666.100 3415.000 2731.900 ;
        RECT 1015.000 2591.900 3415.000 2666.100 ;
        RECT 1015.000 2526.100 1046.390 2591.900 ;
        RECT 1112.040 2526.100 3415.000 2591.900 ;
        RECT 1015.000 2517.900 3415.000 2526.100 ;
        RECT 1015.000 2452.100 3317.960 2517.900 ;
        RECT 3383.610 2452.100 3415.000 2517.900 ;
        RECT 1015.000 2451.900 3415.000 2452.100 ;
        RECT 1015.000 2386.100 1046.390 2451.900 ;
        RECT 1112.040 2386.100 3415.000 2451.900 ;
        RECT 1015.000 2385.900 3415.000 2386.100 ;
        RECT 1015.000 2320.100 3317.960 2385.900 ;
        RECT 3383.610 2320.100 3415.000 2385.900 ;
        RECT 1015.000 2311.900 3415.000 2320.100 ;
        RECT 1015.000 2246.100 1046.390 2311.900 ;
        RECT 1112.040 2253.900 3415.000 2311.900 ;
        RECT 1112.040 2246.100 3317.960 2253.900 ;
        RECT 1015.000 2188.100 3317.960 2246.100 ;
        RECT 3383.610 2188.100 3415.000 2253.900 ;
        RECT 1015.000 2171.900 3415.000 2188.100 ;
        RECT 1015.000 2106.100 1046.390 2171.900 ;
        RECT 1112.040 2121.900 3415.000 2171.900 ;
        RECT 1112.040 2106.100 3317.960 2121.900 ;
        RECT 1015.000 2056.100 3317.960 2106.100 ;
        RECT 3383.610 2056.100 3415.000 2121.900 ;
        RECT 1015.000 2031.900 3415.000 2056.100 ;
        RECT 1015.000 1966.100 1046.390 2031.900 ;
        RECT 1112.040 1989.900 3415.000 2031.900 ;
        RECT 1112.040 1966.100 3317.960 1989.900 ;
        RECT 1015.000 1924.100 3317.960 1966.100 ;
        RECT 3383.610 1924.100 3415.000 1989.900 ;
        RECT 1015.000 1891.900 3415.000 1924.100 ;
        RECT 1015.000 1826.100 1046.390 1891.900 ;
        RECT 1112.040 1857.900 3415.000 1891.900 ;
        RECT 1112.040 1826.100 3317.960 1857.900 ;
        RECT 1015.000 1792.100 3317.960 1826.100 ;
        RECT 3383.610 1792.100 3415.000 1857.900 ;
        RECT 1015.000 1751.900 3415.000 1792.100 ;
        RECT 1015.000 1686.100 1046.390 1751.900 ;
        RECT 1112.040 1725.900 3415.000 1751.900 ;
        RECT 1112.040 1686.100 3317.960 1725.900 ;
        RECT 1015.000 1660.100 3317.960 1686.100 ;
        RECT 3383.610 1660.100 3415.000 1725.900 ;
        RECT 1015.000 1611.900 3415.000 1660.100 ;
        RECT 1015.000 1546.100 1046.390 1611.900 ;
        RECT 1112.040 1593.900 3415.000 1611.900 ;
        RECT 1112.040 1546.100 3317.960 1593.900 ;
        RECT 1015.000 1528.100 3317.960 1546.100 ;
        RECT 3383.610 1528.100 3415.000 1593.900 ;
        RECT 1015.000 1370.090 3415.000 1528.100 ;
        RECT 1015.000 1369.540 2653.600 1370.090 ;
        RECT 1015.000 1303.890 1256.600 1369.540 ;
        RECT 1322.400 1303.890 1373.600 1369.540 ;
        RECT 1439.400 1303.890 1490.600 1369.540 ;
        RECT 1556.400 1303.890 1608.600 1369.540 ;
        RECT 1674.400 1303.890 1725.600 1369.540 ;
        RECT 1791.400 1303.890 1842.600 1369.540 ;
        RECT 1908.400 1303.890 1959.600 1369.540 ;
        RECT 2025.400 1303.890 2077.600 1369.540 ;
        RECT 2143.400 1303.890 2194.600 1369.540 ;
        RECT 2260.400 1303.890 2311.600 1369.540 ;
        RECT 2377.400 1304.275 2653.600 1369.540 ;
        RECT 2719.500 1304.275 3102.600 1370.090 ;
        RECT 3168.500 1304.275 3415.000 1370.090 ;
        RECT 2377.400 1303.890 3415.000 1304.275 ;
        RECT 1015.000 1272.500 3415.000 1303.890 ;
  END
END openram_tc_1kb
END LIBRARY

