VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO hydra
  CLASS BLOCK ;
  FOREIGN hydra ;
  ORIGIN 0.000 0.000 ;
  SIZE 1264.000 BY 1180.000 ;
  PIN DAC_0_VREFL
    PORT
      LAYER MET1 ;
        RECT 176.500 1074.880 229.500 1140.880 ;
    END
  END DAC_0_VREFL
  PIN DAC_0_OUT
    PORT
      LAYER MET1 ;
        RECT 262.500 1074.880 315.500 1140.880 ;
    END
  END DAC_0_OUT
  PIN DAC_0_VREFH
    PORT
      LAYER MET1 ;
        RECT 348.500 1074.880 401.500 1140.880 ;
    END
  END DAC_0_VREFH
  PIN ADC_0_VREFH
    PORT
      LAYER MET1 ;
        RECT 433.500 1074.880 486.500 1140.880 ;
    END
  END ADC_0_VREFH
  PIN ADC_0_IN
    PORT
      LAYER MET1 ;
        RECT 519.500 1074.880 572.500 1140.880 ;
    END
  END ADC_0_IN
  PIN ADC_0_VREFL
    PORT
      LAYER MET1 ;
        RECT 605.500 1074.880 658.500 1140.880 ;
    END
  END ADC_0_VREFL
  PIN DAC_1_VREFL
    PORT
      LAYER MET1 ;
        RECT 776.500 1074.880 829.500 1140.880 ;
    END
  END DAC_1_VREFL
  PIN DAC_1_OUT
    PORT
      LAYER MET1 ;
        RECT 862.500 1074.880 915.500 1140.880 ;
    END
  END DAC_1_OUT
  PIN DAC_1_VREFH
    PORT
      LAYER MET1 ;
        RECT 947.500 1074.880 1000.500 1140.880 ;
    END
  END DAC_1_VREFH
  PIN ADC_1_VREFH
    PORT
      LAYER MET1 ;
        RECT 1158.880 863.500 1224.880 916.500 ;
    END
  END ADC_1_VREFH
  PIN ADC_1_IN
    PORT
      LAYER MET1 ;
        RECT 1158.880 777.500 1224.880 830.500 ;
    END
  END ADC_1_IN
  PIN ADC_1_VREFL
    PORT
      LAYER MET1 ;
        RECT 1158.880 691.500 1224.880 744.500 ;
    END
  END ADC_1_VREFL
  PIN ADC_2_VREFL
    PORT
      LAYER MET1 ;
        RECT 1158.880 434.500 1224.880 487.500 ;
    END
  END ADC_2_VREFL
  PIN ADC_2_IN
    PORT
      LAYER MET1 ;
        RECT 1158.880 348.500 1224.880 401.500 ;
    END
  END ADC_2_IN
  PIN ADC_2_VREFH
    PORT
      LAYER MET1 ;
        RECT 1158.880 262.500 1224.880 315.500 ;
    END
  END ADC_2_VREFH
  PIN DAC_2_VREFH
    PORT
      LAYER MET1 ;
        RECT 947.500 39.120 1000.500 105.120 ;
    END
  END DAC_2_VREFH
  PIN DAC_2_OUT
    PORT
      LAYER MET1 ;
        RECT 862.500 39.120 915.500 105.120 ;
    END
  END DAC_2_OUT
  PIN DAC_2_VREFL
    PORT
      LAYER MET1 ;
        RECT 776.500 39.120 829.500 105.120 ;
    END
  END DAC_2_VREFL
  PIN ADC_3_VREFL
    PORT
      LAYER MET1 ;
        RECT 605.500 39.120 658.500 105.120 ;
    END
  END ADC_3_VREFL
  PIN ADC_3_IN
    PORT
      LAYER MET1 ;
        RECT 519.500 39.120 572.500 105.120 ;
    END
  END ADC_3_IN
  PIN ADC_3_VREFH
    PORT
      LAYER MET1 ;
        RECT 433.500 39.120 486.500 105.120 ;
    END
  END ADC_3_VREFH
  PIN DAC_3_VREFH
    PORT
      LAYER MET1 ;
        RECT 348.500 39.120 401.500 105.120 ;
    END
  END DAC_3_VREFH
  PIN DAC_3_OUT
    PORT
      LAYER MET1 ;
        RECT 262.500 39.120 315.500 105.120 ;
    END
  END DAC_3_OUT
  PIN DAC_3_VREFL
    PORT
      LAYER MET1 ;
        RECT 176.500 39.120 229.500 105.120 ;
    END
  END DAC_3_VREFL
  PIN CSB
    PORT
      LAYER MET1 ;
        RECT 39.120 185.500 105.120 238.500 ;
    END
  END CSB
  PIN SCK
    PORT
      LAYER MET1 ;
        RECT 39.120 279.500 105.120 332.500 ;
    END
  END SCK
  PIN SDI
    PORT
      LAYER MET1 ;
        RECT 39.120 846.500 105.120 899.500 ;
    END
  END SDI
  PIN SDO
    PORT
      LAYER MET1 ;
        RECT 39.120 940.500 105.120 993.500 ;
    END
  END SDO
  PIN VSS
    PORT
      LAYER MET1 ;
        RECT 690.500 1074.880 743.500 1140.880 ;
    END
  END VSS
  PIN VDD1V8
    PORT
      LAYER MET1 ;
        RECT 1033.500 1074.880 1086.500 1140.880 ;
    END
  END VDD1V8
  PIN VDD3V3
    PORT
      LAYER MET1 ;
        RECT 1158.880 949.500 1224.880 1002.500 ;
    END
  END VDD3V3
  OBS
      LAYER MET1 ;
        RECT 0.000 1141.480 1264.000 1180.000 ;
        RECT 0.000 1074.280 175.900 1141.480 ;
        RECT 230.100 1074.280 261.900 1141.480 ;
        RECT 316.100 1074.280 347.900 1141.480 ;
        RECT 402.100 1074.280 432.900 1141.480 ;
        RECT 487.100 1074.280 518.900 1141.480 ;
        RECT 573.100 1074.280 604.900 1141.480 ;
        RECT 659.100 1074.280 689.900 1141.480 ;
        RECT 744.100 1074.280 775.900 1141.480 ;
        RECT 830.100 1074.280 861.900 1141.480 ;
        RECT 916.100 1074.280 946.900 1141.480 ;
        RECT 1001.100 1074.280 1032.900 1141.480 ;
        RECT 1087.100 1074.280 1264.000 1141.480 ;
        RECT 0.000 1003.100 1264.000 1074.280 ;
        RECT 0.000 994.100 1158.280 1003.100 ;
        RECT 0.000 939.900 38.520 994.100 ;
        RECT 105.720 948.900 1158.280 994.100 ;
        RECT 1225.480 948.900 1264.000 1003.100 ;
        RECT 105.720 939.900 1264.000 948.900 ;
        RECT 0.000 917.100 1264.000 939.900 ;
        RECT 0.000 900.100 1158.280 917.100 ;
        RECT 0.000 845.900 38.520 900.100 ;
        RECT 105.720 862.900 1158.280 900.100 ;
        RECT 1225.480 862.900 1264.000 917.100 ;
        RECT 105.720 845.900 1264.000 862.900 ;
        RECT 0.000 831.100 1264.000 845.900 ;
        RECT 0.000 776.900 1158.280 831.100 ;
        RECT 1225.480 776.900 1264.000 831.100 ;
        RECT 0.000 745.100 1264.000 776.900 ;
        RECT 0.000 690.900 1158.280 745.100 ;
        RECT 1225.480 690.900 1264.000 745.100 ;
        RECT 0.000 488.100 1264.000 690.900 ;
        RECT 0.000 433.900 1158.280 488.100 ;
        RECT 1225.480 433.900 1264.000 488.100 ;
        RECT 0.000 402.100 1264.000 433.900 ;
        RECT 0.000 347.900 1158.280 402.100 ;
        RECT 1225.480 347.900 1264.000 402.100 ;
        RECT 0.000 333.100 1264.000 347.900 ;
        RECT 0.000 278.900 38.520 333.100 ;
        RECT 105.720 316.100 1264.000 333.100 ;
        RECT 105.720 278.900 1158.280 316.100 ;
        RECT 0.000 261.900 1158.280 278.900 ;
        RECT 1225.480 261.900 1264.000 316.100 ;
        RECT 0.000 239.100 1264.000 261.900 ;
        RECT 0.000 184.900 38.520 239.100 ;
        RECT 105.720 184.900 1264.000 239.100 ;
        RECT 0.000 105.720 1264.000 184.900 ;
        RECT 0.000 38.520 175.900 105.720 ;
        RECT 230.100 38.520 261.900 105.720 ;
        RECT 316.100 38.520 347.900 105.720 ;
        RECT 402.100 38.520 432.900 105.720 ;
        RECT 487.100 38.520 518.900 105.720 ;
        RECT 573.100 38.520 604.900 105.720 ;
        RECT 659.100 38.520 775.900 105.720 ;
        RECT 830.100 38.520 861.900 105.720 ;
        RECT 916.100 38.520 946.900 105.720 ;
        RECT 1001.100 38.520 1264.000 105.720 ;
        RECT 0.000 0.000 1264.000 38.520 ;
      LAYER MET2 ;
        RECT 0.000 0.000 1264.000 1180.000 ;
      LAYER MET3 ;
        RECT 0.000 0.000 1264.000 1180.000 ;
      LAYER MET4 ;
        RECT 0.000 0.000 1264.000 1180.000 ;
      LAYER METTP ;
        RECT 0.000 0.000 1264.000 1180.000 ;
      LAYER METTPL ;
        RECT 0.000 0.000 1264.000 1180.000 ;
  END
END hydra
END LIBRARY

