VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO striVe2
  CLASS BLOCK ;
  FOREIGN striVe2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2012.000 BY 2041.000 ;
  PIN vdd
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT 225.100 1945.010 287.800 2007.625 ;
    END
  END vdd
  PIN vdd1v8
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT 405.100 1945.010 467.800 2007.625 ;
    END
  END vdd1v8
  PIN vss
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT 495.100 1945.010 557.800 2007.625 ;
    END
  END vss
  PIN gpio[8]
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT 681.200 1945.560 743.800 2008.010 ;
    END
  END gpio[8]
  PIN gpio[7]
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT 776.200 1945.560 838.800 2008.010 ;
    END
  END gpio[7]
  PIN gpio[6]
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT 871.200 1945.560 933.800 2008.010 ;
    END
  END gpio[6]
  PIN gpio[5]
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT 966.200 1945.560 1028.800 2008.010 ;
    END
  END gpio[5]
  PIN gpio[15]
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT 1061.200 1945.560 1123.800 2008.010 ;
    END
  END gpio[15]
  PIN gpio[14]
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT 1156.200 1945.560 1218.800 2008.010 ;
    END
  END gpio[14]
  PIN gpio[13]
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT 1252.200 1945.560 1314.800 2008.010 ;
    END
  END gpio[13]
  PIN gpio[12]
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT 1347.200 1945.560 1409.800 2008.010 ;
    END
  END gpio[12]
  PIN irq
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 1442.200 1945.560 1504.800 2008.010 ;
    END
  END irq
  PIN SDO
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met5 ;
        RECT 1537.200 1945.560 1599.800 2008.010 ;
    END
  END SDO
  PIN SDI
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 1632.200 1945.560 1694.800 2008.010 ;
    END
  END SDI
  PIN flash_csb
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met5 ;
        RECT 1727.200 1945.560 1789.800 2008.010 ;
    END
  END flash_csb
  PIN comp_inn
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 786.200 32.990 848.800 95.440 ;
    END
  END comp_inn
  PIN adc_low
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 900.200 32.990 962.800 95.440 ;
    END
  END adc_low
  PIN adc_high
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 1014.200 32.990 1076.800 95.440 ;
    END
  END adc_high
  PIN adc1_in
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 1128.200 32.990 1190.800 95.440 ;
    END
  END adc1_in
  PIN adc0_in
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 1243.200 32.990 1305.800 95.440 ;
    END
  END adc0_in
  PIN xo
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met5 ;
        RECT 1357.200 32.990 1419.800 95.440 ;
    END
  END xo
  PIN xi
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 1471.200 32.990 1533.800 95.440 ;
    END
  END xi
  PIN gpio[10]
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT 1585.200 32.990 1647.800 95.440 ;
    END
  END gpio[10]
  PIN gpio[9]
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT 1699.200 32.990 1761.800 95.440 ;
    END
  END gpio[9]
  PIN comp_inp
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 32.990 592.200 95.440 654.800 ;
    END
  END comp_inp
  PIN RSTB
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 35.715 693.250 91.545 730.435 ;
    END
  END RSTB
  PIN CSB
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 32.990 777.200 95.440 839.800 ;
    END
  END CSB
  PIN SCK
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 32.990 873.200 95.440 935.800 ;
    END
  END SCK
  PIN xclk
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 32.990 968.200 95.440 1030.800 ;
    END
  END xclk
  PIN flash_clk
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met5 ;
        RECT 32.990 1064.200 95.440 1126.800 ;
    END
  END flash_clk
  PIN flash_io0
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met5 ;
        RECT 32.990 1159.200 95.440 1221.800 ;
    END
  END flash_io0
  PIN flash_io1
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met5 ;
        RECT 32.990 1254.200 95.440 1316.800 ;
    END
  END flash_io1
  PIN flash_io2
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met5 ;
        RECT 32.990 1350.200 95.440 1412.800 ;
    END
  END flash_io2
  PIN flash_io3
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met5 ;
        RECT 32.990 1445.200 95.440 1507.800 ;
    END
  END flash_io3
  PIN ser_rx
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 37.095 1547.930 82.470 1616.325 ;
    END
  END ser_rx
  PIN ser_tx
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met5 ;
        RECT 37.095 1702.930 82.470 1771.325 ;
    END
  END ser_tx
  PIN gpio[4]
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT 1916.560 972.200 1979.010 1034.800 ;
    END
  END gpio[4]
  PIN gpio[3]
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT 1916.560 1117.200 1979.010 1179.800 ;
    END
  END gpio[3]
  PIN gpio[2]
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT 1916.560 1262.200 1979.010 1324.800 ;
    END
  END gpio[2]
  PIN gpio[1]
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT 1916.560 1407.200 1979.010 1469.800 ;
    END
  END gpio[1]
  PIN gpio[0]
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT 1916.560 1552.200 1979.010 1614.800 ;
    END
  END gpio[0]
  PIN gpio[11]
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT 1916.560 1697.200 1979.010 1759.800 ;
    END
  END gpio[11]
  OBS
      LAYER li1 ;
        RECT 0.220 0.220 2011.780 2040.780 ;
      LAYER met1 ;
        RECT 0.000 0.000 2012.000 2041.000 ;
      LAYER met2 ;
        RECT 0.000 0.000 2012.000 2041.000 ;
      LAYER met3 ;
        RECT 0.000 0.000 2012.000 2041.000 ;
      LAYER met4 ;
        RECT 0.000 0.000 2012.000 2041.000 ;
      LAYER met5 ;
        RECT 0.000 2009.610 2012.000 2041.000 ;
        RECT 0.000 2009.225 679.600 2009.610 ;
        RECT 0.000 1943.410 223.500 2009.225 ;
        RECT 289.400 1943.410 403.500 2009.225 ;
        RECT 469.400 1943.410 493.500 2009.225 ;
        RECT 559.400 1943.960 679.600 2009.225 ;
        RECT 745.400 1943.960 774.600 2009.610 ;
        RECT 840.400 1943.960 869.600 2009.610 ;
        RECT 935.400 1943.960 964.600 2009.610 ;
        RECT 1030.400 1943.960 1059.600 2009.610 ;
        RECT 1125.400 1943.960 1154.600 2009.610 ;
        RECT 1220.400 1943.960 1250.600 2009.610 ;
        RECT 1316.400 1943.960 1345.600 2009.610 ;
        RECT 1411.400 1943.960 1440.600 2009.610 ;
        RECT 1506.400 1943.960 1535.600 2009.610 ;
        RECT 1601.400 1943.960 1630.600 2009.610 ;
        RECT 1696.400 1943.960 1725.600 2009.610 ;
        RECT 1791.400 1943.960 2012.000 2009.610 ;
        RECT 559.400 1943.410 2012.000 1943.960 ;
        RECT 0.000 1772.925 2012.000 1943.410 ;
        RECT 0.000 1701.330 35.495 1772.925 ;
        RECT 84.070 1761.400 2012.000 1772.925 ;
        RECT 84.070 1701.330 1914.960 1761.400 ;
        RECT 0.000 1695.600 1914.960 1701.330 ;
        RECT 1980.610 1695.600 2012.000 1761.400 ;
        RECT 0.000 1617.925 2012.000 1695.600 ;
        RECT 0.000 1546.330 35.495 1617.925 ;
        RECT 84.070 1616.400 2012.000 1617.925 ;
        RECT 84.070 1550.600 1914.960 1616.400 ;
        RECT 1980.610 1550.600 2012.000 1616.400 ;
        RECT 84.070 1546.330 2012.000 1550.600 ;
        RECT 0.000 1509.400 2012.000 1546.330 ;
        RECT 0.000 1443.600 31.390 1509.400 ;
        RECT 97.040 1471.400 2012.000 1509.400 ;
        RECT 97.040 1443.600 1914.960 1471.400 ;
        RECT 0.000 1414.400 1914.960 1443.600 ;
        RECT 0.000 1348.600 31.390 1414.400 ;
        RECT 97.040 1405.600 1914.960 1414.400 ;
        RECT 1980.610 1405.600 2012.000 1471.400 ;
        RECT 97.040 1348.600 2012.000 1405.600 ;
        RECT 0.000 1326.400 2012.000 1348.600 ;
        RECT 0.000 1318.400 1914.960 1326.400 ;
        RECT 0.000 1252.600 31.390 1318.400 ;
        RECT 97.040 1260.600 1914.960 1318.400 ;
        RECT 1980.610 1260.600 2012.000 1326.400 ;
        RECT 97.040 1252.600 2012.000 1260.600 ;
        RECT 0.000 1223.400 2012.000 1252.600 ;
        RECT 0.000 1157.600 31.390 1223.400 ;
        RECT 97.040 1181.400 2012.000 1223.400 ;
        RECT 97.040 1157.600 1914.960 1181.400 ;
        RECT 0.000 1128.400 1914.960 1157.600 ;
        RECT 0.000 1062.600 31.390 1128.400 ;
        RECT 97.040 1115.600 1914.960 1128.400 ;
        RECT 1980.610 1115.600 2012.000 1181.400 ;
        RECT 97.040 1062.600 2012.000 1115.600 ;
        RECT 0.000 1036.400 2012.000 1062.600 ;
        RECT 0.000 1032.400 1914.960 1036.400 ;
        RECT 0.000 966.600 31.390 1032.400 ;
        RECT 97.040 970.600 1914.960 1032.400 ;
        RECT 1980.610 970.600 2012.000 1036.400 ;
        RECT 97.040 966.600 2012.000 970.600 ;
        RECT 0.000 937.400 2012.000 966.600 ;
        RECT 0.000 871.600 31.390 937.400 ;
        RECT 97.040 871.600 2012.000 937.400 ;
        RECT 0.000 841.400 2012.000 871.600 ;
        RECT 0.000 775.600 31.390 841.400 ;
        RECT 97.040 775.600 2012.000 841.400 ;
        RECT 0.000 732.035 2012.000 775.600 ;
        RECT 0.000 691.650 34.115 732.035 ;
        RECT 93.145 691.650 2012.000 732.035 ;
        RECT 0.000 656.400 2012.000 691.650 ;
        RECT 0.000 590.600 31.390 656.400 ;
        RECT 97.040 590.600 2012.000 656.400 ;
        RECT 0.000 97.040 2012.000 590.600 ;
        RECT 0.000 31.390 784.600 97.040 ;
        RECT 850.400 31.390 898.600 97.040 ;
        RECT 964.400 31.390 1012.600 97.040 ;
        RECT 1078.400 31.390 1126.600 97.040 ;
        RECT 1192.400 31.390 1241.600 97.040 ;
        RECT 1307.400 31.390 1355.600 97.040 ;
        RECT 1421.400 31.390 1469.600 97.040 ;
        RECT 1535.400 31.390 1583.600 97.040 ;
        RECT 1649.400 31.390 1697.600 97.040 ;
        RECT 1763.400 31.390 2012.000 97.040 ;
        RECT 0.000 0.000 2012.000 31.390 ;
  END
END striVe2
END LIBRARY

