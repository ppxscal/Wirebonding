VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO striVe
  CLASS BLOCK ;
  FOREIGN striVe ;
  ORIGIN 0.000 0.000 ;
  SIZE 2754.000 BY 2762.000 ;
  PIN vdd
    PORT
      LAYER met5 ;
        RECT 39.375 273.100 101.990 335.800 ;
    END
  END vdd
  PIN vss
    PORT
      LAYER met5 ;
        RECT 39.375 669.100 101.990 731.800 ;
    END
  END vss
  PIN comp_inp
    PORT
      LAYER met5 ;
        RECT 38.990 806.200 101.440 868.800 ;
    END
  END comp_inp
  PIN RSTB
    PORT
      LAYER met5 ;
        RECT 41.715 949.250 97.545 986.435 ;
    END
  END RSTB
  PIN CSB
    PORT
      LAYER met5 ;
        RECT 38.990 1075.200 101.440 1137.800 ;
    END
  END CSB
  PIN SCK
    PORT
      LAYER met5 ;
        RECT 38.990 1212.200 101.440 1274.800 ;
    END
  END SCK
  PIN xclk
    PORT
      LAYER met5 ;
        RECT 38.990 1350.200 101.440 1412.800 ;
    END
  END xclk
  PIN flash_clk
    PORT
      LAYER met5 ;
        RECT 38.990 1487.200 101.440 1549.800 ;
    END
  END flash_clk
  PIN flash_io0
    PORT
      LAYER met5 ;
        RECT 38.990 1624.200 101.440 1686.800 ;
    END
  END flash_io0
  PIN flash_io1
    PORT
      LAYER met5 ;
        RECT 38.990 1761.200 101.440 1823.800 ;
    END
  END flash_io1
  PIN flash_io2
    PORT
      LAYER met5 ;
        RECT 38.990 1898.200 101.440 1960.800 ;
    END
  END flash_io2
  PIN flash_io3
    PORT
      LAYER met5 ;
        RECT 38.990 2035.200 101.440 2097.800 ;
    END
  END flash_io3
  PIN ser_rx
    PORT
      LAYER met5 ;
        RECT 43.095 2178.930 88.470 2247.325 ;
    END
  END ser_rx
  PIN ser_tx
    PORT
      LAYER met5 ;
        RECT 43.095 2375.930 88.470 2444.325 ;
    END
  END ser_tx
  PIN gpio[8]
    PORT
      LAYER met5 ;
        RECT 930.200 2660.560 992.800 2723.010 ;
    END
  END gpio[8]
  PIN gpio[7]
    PORT
      LAYER met5 ;
        RECT 1066.200 2660.560 1128.800 2723.010 ;
    END
  END gpio[7]
  PIN gpio[6]
    PORT
      LAYER met5 ;
        RECT 1201.200 2660.560 1263.800 2723.010 ;
    END
  END gpio[6]
  PIN gpio[5]
    PORT
      LAYER met5 ;
        RECT 1337.200 2660.560 1399.800 2723.010 ;
    END
  END gpio[5]
  PIN gpio[15]
    PORT
      LAYER met5 ;
        RECT 1473.200 2660.560 1535.800 2723.010 ;
    END
  END gpio[15]
  PIN gpio[14]
    PORT
      LAYER met5 ;
        RECT 1608.200 2660.560 1670.800 2723.010 ;
    END
  END gpio[14]
  PIN gpio[13]
    PORT
      LAYER met5 ;
        RECT 1744.200 2660.560 1806.800 2723.010 ;
    END
  END gpio[13]
  PIN gpio[12]
    PORT
      LAYER met5 ;
        RECT 1880.200 2660.560 1942.800 2723.010 ;
    END
  END gpio[12]
  PIN irq
    PORT
      LAYER met5 ;
        RECT 2016.200 2660.560 2078.800 2723.010 ;
    END
  END irq
  PIN SDO
    PORT
      LAYER met5 ;
        RECT 2151.200 2660.560 2213.800 2723.010 ;
    END
  END SDO
  PIN SDI
    PORT
      LAYER met5 ;
        RECT 2287.200 2660.560 2349.800 2723.010 ;
    END
  END SDI
  PIN flash_csb
    PORT
      LAYER met5 ;
        RECT 2423.200 2660.560 2485.800 2723.010 ;
    END
  END flash_csb
  PIN gpio[11]
    PORT
      LAYER met5 ;
        RECT 2652.560 2353.200 2715.010 2415.800 ;
    END
  END gpio[11]
  PIN gpio[0]
    PORT
      LAYER met5 ;
        RECT 2652.560 2149.200 2715.010 2211.800 ;
    END
  END gpio[0]
  PIN gpio[1]
    PORT
      LAYER met5 ;
        RECT 2652.560 1945.200 2715.010 2007.800 ;
    END
  END gpio[1]
  PIN gpio[2]
    PORT
      LAYER met5 ;
        RECT 2652.560 1741.200 2715.010 1803.800 ;
    END
  END gpio[2]
  PIN gpio[3]
    PORT
      LAYER met5 ;
        RECT 2652.560 1536.200 2715.010 1598.800 ;
    END
  END gpio[3]
  PIN gpio[4]
    PORT
      LAYER met5 ;
        RECT 2652.560 1332.200 2715.010 1394.800 ;
    END
  END gpio[4]
  PIN gpio[9]
    PORT
      LAYER met5 ;
        RECT 2387.200 38.990 2449.800 101.440 ;
    END
  END gpio[9]
  PIN gpio[10]
    PORT
      LAYER met5 ;
        RECT 2224.200 38.990 2286.800 101.440 ;
    END
  END gpio[10]
  PIN xi
    PORT
      LAYER met5 ;
        RECT 2061.200 38.990 2123.800 101.440 ;
    END
  END xi
  PIN xo
    PORT
      LAYER met5 ;
        RECT 1898.200 38.990 1960.800 101.440 ;
    END
  END xo
  PIN adc0_in
    PORT
      LAYER met5 ;
        RECT 1735.200 38.990 1797.800 101.440 ;
    END
  END adc0_in
  PIN adc1_in
    PORT
      LAYER met5 ;
        RECT 1572.200 38.990 1634.800 101.440 ;
    END
  END adc1_in
  PIN adc_high
    PORT
      LAYER met5 ;
        RECT 1409.200 38.990 1471.800 101.440 ;
    END
  END adc_high
  PIN adc_low
    PORT
      LAYER met5 ;
        RECT 1247.200 38.990 1309.800 101.440 ;
    END
  END adc_low
  PIN comp_inn
    PORT
      LAYER met5 ;
        RECT 1084.200 38.990 1146.800 101.440 ;
    END
  END comp_inn
  PIN vdd1v8
    PORT
      LAYER met5 ;
        RECT 613.045 36.430 669.685 103.860 ;
    END
  END vdd1v8
  OBS
      LAYER li1 ;
        RECT 1.000 1.000 2753.000 2761.000 ;
      LAYER met1 ;
        RECT 1.800 1.800 2752.200 2760.200 ;
      LAYER met2 ;
        RECT 6.000 6.000 2748.000 2756.000 ;
      LAYER met3 ;
        RECT 6.000 6.000 2748.000 2756.000 ;
      LAYER met4 ;
        RECT 6.000 6.000 2748.000 2756.000 ;
      LAYER met5 ;
        RECT 6.000 2724.610 2748.000 2756.000 ;
        RECT 6.000 2658.960 928.600 2724.610 ;
        RECT 994.400 2658.960 1064.600 2724.610 ;
        RECT 1130.400 2658.960 1199.600 2724.610 ;
        RECT 1265.400 2658.960 1335.600 2724.610 ;
        RECT 1401.400 2658.960 1471.600 2724.610 ;
        RECT 1537.400 2658.960 1606.600 2724.610 ;
        RECT 1672.400 2658.960 1742.600 2724.610 ;
        RECT 1808.400 2658.960 1878.600 2724.610 ;
        RECT 1944.400 2658.960 2014.600 2724.610 ;
        RECT 2080.400 2658.960 2149.600 2724.610 ;
        RECT 2215.400 2658.960 2285.600 2724.610 ;
        RECT 2351.400 2658.960 2421.600 2724.610 ;
        RECT 2487.400 2658.960 2748.000 2724.610 ;
        RECT 6.000 2445.925 2748.000 2658.960 ;
        RECT 6.000 2374.330 41.495 2445.925 ;
        RECT 90.070 2417.400 2748.000 2445.925 ;
        RECT 90.070 2374.330 2650.960 2417.400 ;
        RECT 6.000 2351.600 2650.960 2374.330 ;
        RECT 2716.610 2351.600 2748.000 2417.400 ;
        RECT 6.000 2248.925 2748.000 2351.600 ;
        RECT 6.000 2177.330 41.495 2248.925 ;
        RECT 90.070 2213.400 2748.000 2248.925 ;
        RECT 90.070 2177.330 2650.960 2213.400 ;
        RECT 6.000 2147.600 2650.960 2177.330 ;
        RECT 2716.610 2147.600 2748.000 2213.400 ;
        RECT 6.000 2099.400 2748.000 2147.600 ;
        RECT 6.000 2033.600 37.390 2099.400 ;
        RECT 103.040 2033.600 2748.000 2099.400 ;
        RECT 6.000 2009.400 2748.000 2033.600 ;
        RECT 6.000 1962.400 2650.960 2009.400 ;
        RECT 6.000 1896.600 37.390 1962.400 ;
        RECT 103.040 1943.600 2650.960 1962.400 ;
        RECT 2716.610 1943.600 2748.000 2009.400 ;
        RECT 103.040 1896.600 2748.000 1943.600 ;
        RECT 6.000 1825.400 2748.000 1896.600 ;
        RECT 6.000 1759.600 37.390 1825.400 ;
        RECT 103.040 1805.400 2748.000 1825.400 ;
        RECT 103.040 1759.600 2650.960 1805.400 ;
        RECT 6.000 1739.600 2650.960 1759.600 ;
        RECT 2716.610 1739.600 2748.000 1805.400 ;
        RECT 6.000 1688.400 2748.000 1739.600 ;
        RECT 6.000 1622.600 37.390 1688.400 ;
        RECT 103.040 1622.600 2748.000 1688.400 ;
        RECT 6.000 1600.400 2748.000 1622.600 ;
        RECT 6.000 1551.400 2650.960 1600.400 ;
        RECT 6.000 1485.600 37.390 1551.400 ;
        RECT 103.040 1534.600 2650.960 1551.400 ;
        RECT 2716.610 1534.600 2748.000 1600.400 ;
        RECT 103.040 1485.600 2748.000 1534.600 ;
        RECT 6.000 1414.400 2748.000 1485.600 ;
        RECT 6.000 1348.600 37.390 1414.400 ;
        RECT 103.040 1396.400 2748.000 1414.400 ;
        RECT 103.040 1348.600 2650.960 1396.400 ;
        RECT 6.000 1330.600 2650.960 1348.600 ;
        RECT 2716.610 1330.600 2748.000 1396.400 ;
        RECT 6.000 1276.400 2748.000 1330.600 ;
        RECT 6.000 1210.600 37.390 1276.400 ;
        RECT 103.040 1210.600 2748.000 1276.400 ;
        RECT 6.000 1139.400 2748.000 1210.600 ;
        RECT 6.000 1073.600 37.390 1139.400 ;
        RECT 103.040 1073.600 2748.000 1139.400 ;
        RECT 6.000 988.035 2748.000 1073.600 ;
        RECT 6.000 947.650 40.115 988.035 ;
        RECT 99.145 947.650 2748.000 988.035 ;
        RECT 6.000 870.400 2748.000 947.650 ;
        RECT 6.000 804.600 37.390 870.400 ;
        RECT 103.040 804.600 2748.000 870.400 ;
        RECT 6.000 733.400 2748.000 804.600 ;
        RECT 6.000 667.500 37.775 733.400 ;
        RECT 103.590 667.500 2748.000 733.400 ;
        RECT 6.000 337.400 2748.000 667.500 ;
        RECT 6.000 271.500 37.775 337.400 ;
        RECT 103.590 271.500 2748.000 337.400 ;
        RECT 6.000 105.460 2748.000 271.500 ;
        RECT 6.000 34.830 611.445 105.460 ;
        RECT 671.285 103.040 2748.000 105.460 ;
        RECT 671.285 37.390 1082.600 103.040 ;
        RECT 1148.400 37.390 1245.600 103.040 ;
        RECT 1311.400 37.390 1407.600 103.040 ;
        RECT 1473.400 37.390 1570.600 103.040 ;
        RECT 1636.400 37.390 1733.600 103.040 ;
        RECT 1799.400 37.390 1896.600 103.040 ;
        RECT 1962.400 37.390 2059.600 103.040 ;
        RECT 2125.400 37.390 2222.600 103.040 ;
        RECT 2288.400 37.390 2385.600 103.040 ;
        RECT 2451.400 37.390 2748.000 103.040 ;
        RECT 671.285 34.830 2748.000 37.390 ;
        RECT 6.000 6.000 2748.000 34.830 ;
  END
END striVe
END LIBRARY

